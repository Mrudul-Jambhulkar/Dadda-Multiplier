module dadda(
input [15:0] a, 
input [15:0] b, 
 output [31:0] y 
);



wire [15:0] pp [0:15];
genvar j ;

for(j=0;j<16;j=j+1)
begin:loop1
assign pp[j][15:0] = ( { 16{b[j]} } & a[15:0] );
end

assign p = pp[14];

wire  c0_0 ; wire [1:0] c0_1 ; wire [2:0] c0_2 ; wire [3:0] c0_3 ; wire [4:0] c0_4 ; wire [5:0] c0_5 ; wire [6:0] c0_6 ; wire [7:0] c0_7 ;

wire [8:0] c0_8 ; wire [9:0] c0_9 ; wire [10:0] c0_10 ; wire [11:0] c0_11;  wire [12:0] c0_12 ; wire [13:0] c0_13 ; wire [14:0] c0_14 ; wire [15:0] c0_15 ;

wire [15:1] c0_16 ; wire [15:2] c0_17 ;  wire [15:3] c0_18 ; wire [15:4] c0_19 ; wire [15:5] c0_20 ; wire [15:6] c0_21 ; wire [15:7] c0_22 ; wire [15:8] c0_23 ; 

wire [15:9] c0_24 ; wire [15:10] c0_25 ;  wire [15:11] c0_26 ; wire [15:12] c0_27 ; wire [15:13] c0_28 ; wire [15:14] c0_29 ; wire  c0_30 ; 

assign c0_0 = pp[0][0];
assign c0_1[1:0] = {pp[0][1],pp[1][0]};
assign c0_2[2:0] = {pp[0][2],pp[1][1],pp[2][0]};
assign c0_3[3:0] = {pp[0][3],pp[1][2],pp[2][1],pp[3][0]};
assign c0_4[4:0] = {pp[0][4],pp[1][3],pp[2][2],pp[3][1],pp[4][0]};
assign c0_5[5:0] = {pp[0][5],pp[1][4],pp[2][3],pp[3][2],pp[4][1],pp[5][0]};
assign c0_6[6:0] = {pp[0][6],pp[1][5],pp[2][4],pp[3][3],pp[4][2],pp[5][1],pp[6][0]};
assign c0_7[7:0] = {pp[0][7],pp[1][6],pp[2][5],pp[3][4],pp[4][3],pp[5][2],pp[6][1],pp[7][0]};
assign c0_8[8:0] = {pp[0][8],pp[1][7],pp[2][6],pp[3][5],pp[4][4],pp[5][3],pp[6][2],pp[7][1],pp[8][0]};
assign c0_9[9:0] = {pp[0][9],pp[1][8],pp[2][7],pp[3][6],pp[4][5],pp[5][4],pp[6][3],pp[7][2],pp[8][1],pp[9][0]};
assign c0_10[10:0] = {pp[0][10],pp[1][9],pp[2][8],pp[3][7],pp[4][6],pp[5][5],pp[6][4],pp[7][3],pp[8][2],pp[9][1],pp[10][0]};
assign c0_11[11:0] = {pp[0][11],pp[1][10],pp[2][9],pp[3][8],pp[4][7],pp[5][6],pp[6][5],pp[7][4],pp[8][3],pp[9][2],pp[10][1],pp[11][0]};
assign c0_12[12:0] = {pp[0][12],pp[1][11],pp[2][10],pp[3][9],pp[4][8],pp[5][7],pp[6][6],pp[7][5],pp[8][4],pp[9][3],pp[10][2],pp[11][1],pp[12][0]};
assign c0_13[13:0] = {pp[0][13],pp[1][12],pp[2][11],pp[3][10],pp[4][9],pp[5][8],pp[6][7],pp[7][6],pp[8][5],pp[9][4],pp[10][3],pp[11][2],pp[12][1],pp[13][0]};
assign c0_14[14:0] = {pp[0][14],pp[1][13],pp[2][12],pp[3][11],pp[4][10],pp[5][9],pp[6][8],pp[7][7],pp[8][6],pp[9][5],pp[10][4],pp[11][3],pp[12][2],pp[13][1],pp[14][0]};
assign c0_15[15:0] = {pp[0][15],pp[1][14],pp[2][13],pp[3][12],pp[4][11],pp[5][10],pp[6][9],pp[7][8],pp[8][7],pp[9][6],pp[10][5],pp[11][4],pp[12][3],pp[13][2],pp[14][1],pp[15][0]};

assign c0_16[15:1] = {pp[1][15],pp[2][14],pp[3][13],pp[4][12],pp[5][11],pp[6][10],pp[7][9],pp[8][8],pp[9][7],pp[10][6],pp[11][5],pp[12][4],pp[13][3],pp[14][2],pp[15][1]};
assign c0_17[15:2] = {pp[2][15],pp[3][14],pp[4][13],pp[5][12],pp[6][11],pp[7][10],pp[8][9],pp[9][8],pp[10][7],pp[11][6],pp[12][5],pp[13][4],pp[14][3],pp[15][2]};
assign c0_18[15:3] = {pp[3][15],pp[4][14],pp[5][13],pp[6][12],pp[7][11],pp[8][10],pp[9][9],pp[10][8],pp[11][7],pp[12][6],pp[13][5],pp[14][4],pp[15][3]};
assign c0_19[15:4] = {pp[4][15],pp[5][14],pp[6][13],pp[7][12],pp[8][11],pp[9][10],pp[10][9],pp[11][8],pp[12][7],pp[13][6],pp[14][5],pp[15][4]};
assign c0_20[15:5] = {pp[5][15],pp[6][14],pp[7][13],pp[8][12],pp[9][11],pp[10][10],pp[11][9],pp[12][8],pp[13][7],pp[14][6],pp[15][5]};
assign c0_21[15:6] = {pp[6][15],pp[7][14],pp[8][13],pp[9][12],pp[10][11],pp[11][10],pp[12][9],pp[13][8],pp[14][7],pp[15][6]};
assign c0_22[15:7] = {pp[7][15],pp[8][14],pp[9][13],pp[10][12],pp[11][11],pp[12][10],pp[13][9],pp[14][8],pp[15][7]};
assign c0_23[15:8] = {pp[8][15],pp[9][14],pp[10][13],pp[11][12],pp[12][11],pp[13][10],pp[14][9],pp[15][8]};
assign c0_24[15:9] = {pp[9][15],pp[10][14],pp[11][13],pp[12][12],pp[13][11],pp[14][10],pp[15][9]};
assign c0_25[15:10] = {pp[10][15],pp[11][14],pp[12][13],pp[13][12],pp[14][11],pp[15][10]};
assign c0_26[15:11] = {pp[11][15],pp[12][14],pp[13][13],pp[14][12],pp[15][11]};
assign c0_27[15:12] = {pp[12][15],pp[13][14],pp[14][13],pp[15][12]};
assign c0_28[15:13] = {pp[13][15],pp[14][14],pp[15][13]};
assign c0_29[15:14] = {pp[14][15],pp[15][14]};
assign c0_30= pp[15][15];


//STAGE 1
wire  c1_0 ; wire [1:0] c1_1 ; wire [2:0] c1_2 ; wire [3:0] c1_3 ; wire [4:0] c1_4 ; wire [5:0] c1_5 ; wire [6:0] c1_6 ; wire [7:0] c1_7 ;

wire [8:0] c1_8 ; wire [9:0] c1_9 ; wire [10:0] c1_10 ; wire [11:0] c1_11;  wire [12:1] c1_12 ; wire [13:2] c1_13 ; wire [14:3] c1_14 ; wire [15:4] c1_15 ;

wire [16:5] c1_16 ; wire [17:6] c1_17 ;  wire [18:7] c1_18 ; wire [19:8] c1_19 ; wire [20:9] c1_20 ; wire [21:12] c1_21 ; wire [22:14] c1_22 ; wire [23:16] c1_23 ; 

wire [24:18] c1_24 ; wire [25:20] c1_25 ;  wire [26:22] c1_26 ; wire [27:24] c1_27 ; wire [28:26] c1_28 ; wire [29:28] c1_29 ; wire  c1_30 ; 

assign c1_0=c0_0 ; assign c1_1=c0_1 ; assign c1_2 = c0_2 ; assign c1_3 = c0_3 ; assign c1_4 = c0_4 ; assign c1_5=c0_5; assign c1_6 = c0_6 ; assign c1_7=c0_7 ;assign c1_8=c0_8;
assign c1_9=c0_9; assign c1_10=c0_10; assign c1_11=c0_11 ;

//idx 12
halfAdder ha1 (.a(c0_12[12]) , .b(c0_12[11]) , .s(c1_12[12]) , .c(c1_13[13]) ) ;
assign c1_12[11:1]=c0_12[10:0];

//idx 13
fullAdder fa1 (.a(c0_13[13]) , .b(c0_13[12]) , .cin(c0_13[11]) , .s(c1_13[12]) , .c(c1_14[14]) ) ;
halfAdder ha2 (.a(c0_13[10]) , .b(c0_13[9]) , .s(c1_13[11]) , .c(c1_14[13]) ) ;
assign c1_13[10:2] = c0_13[8:0];

//idx 14
fullAdder fa2 (.a(c0_14[14]) , .b(c0_14[13]) , .cin(c0_14[12]) , .s(c1_14[12]) , .c(c1_15[15]) ) ;
fullAdder fa3 (.a(c0_14[11]) , .b(c0_14[10]) , .cin(c0_14[9]) , .s(c1_14[11]) , .c(c1_15[14]) ) ;
halfAdder ha3 (.a(c0_14[8]) , .b(c0_14[7]) , .s(c1_14[10]) , .c(c1_15[13]) ) ;
assign c1_14[9:3]=c0_14[6:0];

//idx 15
fullAdder fa4 (.a(c0_15[15]) , .b(c0_15[14]) , .cin(c0_15[13]) , .s(c1_15[12]) , .c(c1_16[16]) ) ;
fullAdder fa5 (.a(c0_15[12]) , .b(c0_15[11]) , .cin(c0_15[10]) , .s(c1_15[11]) , .c(c1_16[15]) ) ;
fullAdder fa6 (.a(c0_15[9]) , .b(c0_15[8]) , .cin(c0_15[7]) , .s(c1_15[10]) , .c(c1_16[14]) ) ;
halfAdder ha4 (.a(c0_15[6]) , .b(c0_15[5]) , .s(c1_15[9]) , .c(c1_16[13]) ) ;
assign c1_15[8:4] = c0_15[4:0];

//idx 16
fullAdder fa7 (.a(c0_16[15]) , .b(c0_16[14]) , .cin(c0_16[13]) , .s(c1_16[12]) , .c(c1_17[17]) ) ;
fullAdder fa8 (.a(c0_16[12]) , .b(c0_16[11]) , .cin(c0_16[10]) , .s(c1_16[11]) , .c(c1_17[16]) ) ;
fullAdder fa9 (.a(c0_16[9]) , .b(c0_16[8]) , .cin(c0_16[7]) , .s(c1_16[10]) , .c(c1_17[15]) ) ;
halfAdder ha5 (.a(c0_16[6]) , .b(c0_16[5]) , .s(c1_16[9]) , .c(c1_17[14]) ) ;
assign c1_16[8:5] = c0_16[4:1];

//idx 17
fullAdder fa10 (.a(c0_17[15]) , .b(c0_17[14]) , .cin(c0_17[13]) , .s(c1_17[13]) , .c(c1_18[18]) ) ;
fullAdder fa11 (.a(c0_17[12]) , .b(c0_17[11]) , .cin(c0_17[10]) , .s(c1_17[12]) , .c(c1_18[17]) ) ;
fullAdder fa12 (.a(c0_17[9]) , .b(c0_17[8]) , .cin(c0_17[7]) , .s(c1_17[11]) , .c(c1_18[16]) ) ;
assign c1_17[10:6] = c0_17[6:2];

//idx 18
fullAdder fa13 (.a(c0_18[15]) , .b(c0_18[14]) , .cin(c0_18[13]) , .s(c1_18[15]) , .c(c1_19[19]) ) ;
fullAdder fa14 (.a(c0_18[12]) , .b(c0_18[11]) , .cin(c0_18[10]) , .s(c1_18[14]) , .c(c1_19[18]) ) ;
assign c1_18[13:7] = c0_18[9:3];

//idx 19
fullAdder fa15 (.a(c0_19[15]) , .b(c0_19[14]) , .cin(c0_19[13]) , .s(c1_19[17]) , .c(c1_20[20]) ) ;
assign c1_19[16:8]=c0_19[12:4] ;

assign c1_20[19:9]=c0_20[15:5];
assign c1_21[21:12]=c0_21[15:6];
assign c1_22[22:14]=c0_22[15:7];
assign c1_23[23:16]=c0_23[15:8];
assign c1_24[24:18]=c0_24[15:9];
assign c1_25[25:20]=c0_25[15:10];
assign c1_26[26:22]=c0_26[15:11];

assign c1_27[27:24]=c0_27[15:12];
assign c1_28[28:26]=c0_28[15:13];
assign c1_29[29:28]=c0_29[15:14];
assign c1_30 = c0_30;




//STAGE 2
wire  c2_0 ; wire [1:0] c2_1 ; wire [2:0] c2_2 ; wire [3:0] c2_3 ; wire [4:0] c2_4 ; wire [5:0] c2_5 ; wire [6:0] c2_6 ; wire [7:0] c2_7 ;

wire [8:0] c2_8 ; wire [9:1] c2_9 ; wire [10:2] c2_10 ; wire [11:3] c2_11;  wire [12:4] c2_12 ; wire [13:5] c2_13 ; wire [14:6] c2_14 ; wire [15:7] c2_15 ;

wire [16:8] c2_16 ; wire [17:9] c2_17 ;  wire [18:10] c2_18 ; wire [19:11] c2_19 ; wire [20:12] c2_20 ; wire [21:13] c2_21 ; wire [22:14] c2_22 ; wire [23:15] c2_23; 

wire [24:18] c2_24 ; wire [25:20] c2_25 ;  wire [26:22] c2_26 ; wire [27:24] c2_27 ; wire [28:26] c2_28 ; wire [29:28] c2_29 ; wire  c2_30 ; 

assign c2_0=c1_0 ; assign c2_1=c1_1 ; assign c2_2 = c1_2 ; assign c2_3 = c1_3 ; assign c2_4 = c1_4 ; assign c2_5=c1_5; assign c2_6 = c1_6 ; assign c2_7=c1_7 ;assign c2_8=c1_8;

//idx9
halfAdder ha2_1 (.a(c1_9[9]) , .b(c1_9[8]) , .s(c2_9[9]) , .c(c2_10[10]) ) ;
assign c2_9[8:1]=c1_9[7:0];

//idx 10
fullAdder fa2_1 (.a(c1_10[10]) , .b(c1_10[9]) , .cin(c1_10[8]) , .s(c2_10[9]) , .c(c2_11[11]) ) ;
halfAdder ha2_2 (.a(c1_10[7]) , .b(c1_10[6]) , .s(c2_10[8]) , .c(c2_11[10]) ) ;
assign c2_10[7:2] = c1_10[5:0];

//idx 11
fullAdder fa2_2 (.a(c1_11[11]) , .b(c1_11[10]) , .cin(c1_11[9]) , .s(c2_11[9]) , .c(c2_12[12]) ) ;
fullAdder fa2_3 (.a(c1_11[8]) , .b(c1_11[7]) , .cin(c1_11[6]) , .s(c2_11[8]) , .c(c2_12[11]) ) ;
halfAdder ha2_3 (.a(c1_11[5]) , .b(c1_11[4]) , .s(c2_11[7]) , .c(c2_12[10]) ) ;
assign c2_11[6:3] = c1_11[3:0];

//idx 12
fullAdder fa2_4 (.a(c1_12[12]) , .b(c1_12[11]) , .cin(c1_12[10]) , .s(c2_12[9]) , .c(c2_13[13]) ) ;
fullAdder fa2_5 (.a(c1_12[9]) , .b(c1_12[8]) , .cin(c1_12[7]) , .s(c2_12[8]) , .c(c2_13[12]) ) ;
fullAdder fa2_6 (.a(c1_12[6]) , .b(c1_12[5]) , .cin(c1_12[4]) , .s(c2_12[7]) , .c(c2_13[11]) ) ;
assign c2_12[6:4] = c1_12[3:1];

//idx 13
fullAdder fa2_7 (.a(c1_13[13]) , .b(c1_13[12]) , .cin(c1_13[11]) , .s(c2_13[10]) , .c(c2_14[14]) ) ;
fullAdder fa2_8 (.a(c1_13[10]) , .b(c1_13[9]) , .cin(c1_13[8]) , .s(c2_13[9]) , .c(c2_14[13]) ) ;
fullAdder fa2_9 (.a(c1_13[7]) , .b(c1_13[6]) , .cin(c1_13[5]) , .s(c2_13[8]) , .c(c2_14[12]) ) ;
assign c2_13[7:5] = c1_13[4:2];

//idx 14
fullAdder fa2_10 (.a(c1_14[14]) , .b(c1_14[13]) , .cin(c1_14[12]) , .s(c2_14[11]) , .c(c2_15[15]) ) ;
fullAdder fa2_11 (.a(c1_14[11]) , .b(c1_14[10]) , .cin(c1_14[9]) , .s(c2_14[10]) , .c(c2_15[14]) ) ;
fullAdder fa2_12 (.a(c1_14[8]) , .b(c1_14[7]) , .cin(c1_14[6]) , .s(c2_14[9]) , .c(c2_15[13]) ) ;
assign c2_14[8:6] = c1_14[5:3];

//idx 15
fullAdder fa2_13 (.a(c1_15[15]) , .b(c1_15[14]) , .cin(c1_15[13]) , .s(c2_15[12]) , .c(c2_16[16]) ) ;
fullAdder fa2_14 (.a(c1_15[12]) , .b(c1_15[11]) , .cin(c1_15[10]) , .s(c2_15[11]) , .c(c2_16[15]) ) ;
fullAdder fa2_15 (.a(c1_15[9]) , .b(c1_15[8]) , .cin(c1_15[7]) , .s(c2_15[10]) , .c(c2_16[14]) ) ;
assign c2_15[9:7] = c1_15[6:4];

//idx 16
fullAdder fa2_16 (.a(c1_16[16]) , .b(c1_16[15]) , .cin(c1_16[14]) , .s(c2_16[13]) , .c(c2_17[17]) ) ;
fullAdder fa2_17 (.a(c1_16[13]) , .b(c1_16[12]) , .cin(c1_16[11]) , .s(c2_16[12]) , .c(c2_17[16]) ) ;
fullAdder fa2_18 (.a(c1_16[10]) , .b(c1_16[9]) , .cin(c1_16[8]) , .s(c2_16[11]) , .c(c2_17[15]) ) ;
assign c2_16[10:8] = c1_16[7:5];

//idx 17
fullAdder fa2_19 (.a(c1_17[17]) , .b(c1_17[16]) , .cin(c1_17[15]) , .s(c2_17[14]) , .c(c2_18[18]) ) ;
fullAdder fa2_20 (.a(c1_17[14]) , .b(c1_17[13]) , .cin(c1_17[12]) , .s(c2_17[13]) , .c(c2_18[17]) ) ;
fullAdder fa2_21 (.a(c1_17[11]) , .b(c1_17[10]) , .cin(c1_17[9]) , .s(c2_17[12]) , .c(c2_18[16]) ) ;
assign c2_17[11:9] = c1_17[8:6];

//idx 18
fullAdder fa2_22 (.a(c1_18[18]) , .b(c1_18[17]) , .cin(c1_18[16]) , .s(c2_18[15]) , .c(c2_19[19]) ) ;
fullAdder fa2_23 (.a(c1_18[15]) , .b(c1_18[14]) , .cin(c1_18[13]) , .s(c2_18[14]) , .c(c2_19[18]) ) ;
fullAdder fa2_24 (.a(c1_18[12]) , .b(c1_18[11]) , .cin(c1_18[10]) , .s(c2_18[13]) , .c(c2_19[17]) ) ;
assign c2_18[12:10] = c1_18[9:7];

//idx 19
fullAdder fa2_25 (.a(c1_19[19]) , .b(c1_19[18]) , .cin(c1_19[17]) , .s(c2_19[16]) , .c(c2_20[20]) ) ;
fullAdder fa2_26 (.a(c1_19[16]) , .b(c1_19[15]) , .cin(c1_19[14]) , .s(c2_19[15]) , .c(c2_20[19]) ) ;
fullAdder fa2_27 (.a(c1_19[13]) , .b(c1_19[12]) , .cin(c1_19[11]) , .s(c2_19[14]) , .c(c2_20[18]) ) ;
assign c2_19[13:11] = c1_19[10:8];

//idx 20
fullAdder fa2_28 (.a(c1_20[20]) , .b(c1_20[19]) , .cin(c1_20[18]) , .s(c2_20[17]) , .c(c2_21[21]) ) ;
fullAdder fa2_29 (.a(c1_20[17]) , .b(c1_20[16]) , .cin(c1_20[15]) , .s(c2_20[16]) , .c(c2_21[20]) ) ;
fullAdder fa2_30 (.a(c1_20[14]) , .b(c1_20[13]) , .cin(c1_20[12]) , .s(c2_20[15]) , .c(c2_21[19]) ) ;
assign c2_20[14:12] = c1_20[11:9];

//idx 21
fullAdder fa2_31 (.a(c1_21[21]) , .b(c1_21[20]) , .cin(c1_21[19]) , .s(c2_21[18]) , .c(c2_22[22]) ) ;
fullAdder fa2_32 (.a(c1_21[18]) , .b(c1_21[17]) , .cin(c1_21[16]) , .s(c2_21[17]) , .c(c2_22[21]) ) ;
assign c2_21[16:13]=c1_21[15:12] ;

//idx 22
fullAdder fa2_33 (.a(c1_22[22]) , .b(c1_22[21]) , .cin(c1_22[20]) , .s(c2_22[20]) , .c(c2_23[23]) ) ;
assign c2_22[19:14]=c1_22[19:14] ;

//idx 23
assign c2_23[22:15]=c1_23[23:16];

assign c2_24[24:18]=c1_24[24:18];
assign c2_25[25:20]=c1_25[25:20];
assign c2_26[26:22]=c1_26[26:22];
assign c2_27[27:24]=c1_27[27:24];
assign c2_28[28:26]=c1_28[28:26];
assign c2_29[29:28]=c1_29[29:28];
assign c2_30 = c1_30 ;

//STAGE 3
wire  c3_0 ; wire [1:0] c3_1 ; wire [2:0] c3_2 ; wire [3:0] c3_3 ; wire [4:0] c3_4 ; wire [5:0] c3_5 ; wire [6:1] c3_6 ; wire [7:2] c3_7 ;

wire [8:3] c3_8 ; wire [9:4] c3_9 ; wire [10:5] c3_10 ; wire [11:6] c3_11;  wire [12:7] c3_12 ; wire [13:8] c3_13 ; wire [14:9] c3_14 ; wire [15:10] c3_15 ;

wire [16:11] c3_16; wire [17:12] c3_17; wire [18:13] c3_18; wire [19:14] c3_19; wire [20:15] c3_20; wire [21:16] c3_21; wire [22:17] c3_22; wire [23:18] c3_23; 
wire [24:19] c3_24; wire [25:20] c3_25; wire [26:21] c3_26; wire [27:24] c3_27 ; wire [28:26] c3_28 ; wire [29:28] c3_29 ; wire  c3_30 ;

assign c3_0 = c2_0 ; assign c3_1 = c2_1; assign c3_2 = c2_2 ; assign c3_3 = c2_3; assign c3_4 = c2_4 ; assign c3_5 = c2_5;

//idx6
halfAdder ha3_1 (.a(c2_6[6]) , .b(c2_6[5]) , .s(c3_6[6]) , .c(c3_7[7]) ) ;
assign c3_6[5:1]=c2_6[4:0];

//idx7
fullAdder fa3_1 (.a(c2_7[7]) , .b(c2_7[6]) , .cin(c2_7[5]) , .s(c3_7[6]) , .c(c3_8[8]) ) ;
halfAdder ha3_2 (.a(c2_7[4]) , .b(c2_7[3]) , .s(c3_7[5]) , .c(c3_8[7]) ) ;
assign c3_7[4:2] = c2_7[2:0];

//idx8
fullAdder fa3_2 (.a(c2_8[8]) , .b(c2_8[7]) , .cin(c2_8[6]) , .s(c3_8[6]) , .c(c3_9[9]) ) ;
fullAdder fa3_3 (.a(c2_8[5]) , .b(c2_8[4]) , .cin(c2_8[3]) , .s(c3_8[5]) , .c(c3_9[8]) ) ;
halfAdder ha3_3 (.a(c2_8[2]) , .b(c2_8[1]) , .s(c3_8[4]) , .c(c3_9[7]) ) ;
assign c3_8[3] = c2_8[0];

//idx9
fullAdder fa3_4 (.a(c2_9[9]) , .b(c2_9[8]) , .cin(c2_9[7]) , .s(c3_9[6]) , .c(c3_10[10]) ) ;
fullAdder fa3_5 (.a(c2_9[6]) , .b(c2_9[5]) , .cin(c2_9[4]) , .s(c3_9[5]) , .c(c3_10[9]) ) ;
fullAdder fa3_6 (.a(c2_9[3]) , .b(c2_9[2]) , .cin(c2_9[1]) , .s(c3_9[4]) , .c(c3_10[8]) ) ;

//idx10
fullAdder fa3_7 (.a(c2_10[10]) , .b(c2_10[9]) , .cin(c2_10[8]) , .s(c3_10[7]) , .c(c3_11[11]) ) ;
fullAdder fa3_8 (.a(c2_10[7]) , .b(c2_10[6]) , .cin(c2_10[5]) , .s(c3_10[6]) , .c(c3_11[10]) ) ;
fullAdder fa3_9 (.a(c2_10[4]) , .b(c2_10[3]) , .cin(c2_10[2]) , .s(c3_10[5]) , .c(c3_11[9]) ) ;

//continue
//idx11
fullAdder fa3_10 (.a(c2_11[11]) , .b(c2_11[10]) , .cin(c2_11[9]) , .s(c3_11[8]) , .c(c3_12[12]) ) ;
fullAdder fa3_11 (.a(c2_11[8]) , .b(c2_11[7]) , .cin(c2_11[6]) , .s(c3_11[7]) , .c(c3_12[11]) ) ;
fullAdder fa3_12 (.a(c2_11[5]) , .b(c2_11[4]) , .cin(c2_11[3]) , .s(c3_11[6]) , .c(c3_12[10]) ) ;

//idx12
fullAdder fa3_13 (.a(c2_12[12]) , .b(c2_12[11]) , .cin(c2_12[10]) , .s(c3_12[9]) , .c(c3_13[13]) ) ;
fullAdder fa3_14 (.a(c2_12[9]) , .b(c2_12[8]) , .cin(c2_12[7]) , .s(c3_12[8]) , .c(c3_13[12]) ) ;
fullAdder fa3_15 (.a(c2_12[6]) , .b(c2_12[5]) , .cin(c2_12[4]) , .s(c3_12[7]) , .c(c3_13[11]) ) ;

//idx13
fullAdder fa3_16 (.a(c2_13[13]) , .b(c2_13[12]) , .cin(c2_13[11]) , .s(c3_13[10]) , .c(c3_14[14]) ) ;
fullAdder fa3_17 (.a(c2_13[10]) , .b(c2_13[9]) , .cin(c2_13[8]) , .s(c3_13[9]) , .c(c3_14[13]) ) ;
fullAdder fa3_18 (.a(c2_13[7]) , .b(c2_13[6]) , .cin(c2_13[5]) , .s(c3_13[8]) , .c(c3_14[12]) ) ;

//idx14
fullAdder fa3_19 (.a(c2_14[14]) , .b(c2_14[13]) , .cin(c2_14[12]) , .s(c3_14[11]) , .c(c3_15[15]) ) ;
fullAdder fa3_20 (.a(c2_14[11]) , .b(c2_14[10]) , .cin(c2_14[9]) , .s(c3_14[10]) , .c(c3_15[14]) ) ;
fullAdder fa3_21 (.a(c2_14[8]) , .b(c2_14[7]) , .cin(c2_14[6]) , .s(c3_14[9]) , .c(c3_15[13]) ) ;

//idx15
fullAdder fa3_22 (.a(c2_15[15]) , .b(c2_15[14]) , .cin(c2_15[13]) , .s(c3_15[12]) , .c(c3_16[16]) ) ;
fullAdder fa3_23 (.a(c2_15[12]) , .b(c2_15[11]) , .cin(c2_15[10]) , .s(c3_15[11]) , .c(c3_16[15]) ) ;
fullAdder fa3_24 (.a(c2_15[9]) , .b(c2_15[8]) , .cin(c2_15[7]) , .s(c3_15[10]) , .c(c3_16[14]) ) ;

//idx16
fullAdder fa3_25 (.a(c2_16[16]) , .b(c2_16[15]) , .cin(c2_16[14]) , .s(c3_16[13]) , .c(c3_17[17]) ) ;
fullAdder fa3_26 (.a(c2_16[13]) , .b(c2_16[12]) , .cin(c2_16[11]) , .s(c3_16[12]) , .c(c3_17[16]) ) ;
fullAdder fa3_27 (.a(c2_16[10]) , .b(c2_16[9]) , .cin(c2_16[8]) , .s(c3_16[11]) , .c(c3_17[15]) ) ;

//idx17
fullAdder fa3_28 (.a(c2_17[17]) , .b(c2_17[16]) , .cin(c2_17[15]) , .s(c3_17[14]) , .c(c3_18[18]) ) ;
fullAdder fa3_29 (.a(c2_17[14]) , .b(c2_17[13]) , .cin(c2_17[12]) , .s(c3_17[13]) , .c(c3_18[17]) ) ;
fullAdder fa3_30 (.a(c2_17[11]) , .b(c2_17[10]) , .cin(c2_17[9]) , .s(c3_17[12]) , .c(c3_18[16]) ) ;

//idx18
fullAdder fa3_31 (.a(c2_18[18]) , .b(c2_18[17]) , .cin(c2_18[16]) , .s(c3_18[15]) , .c(c3_19[19]) ) ;
fullAdder fa3_32 (.a(c2_18[15]) , .b(c2_18[14]) , .cin(c2_18[13]) , .s(c3_18[14]) , .c(c3_19[18]) ) ;
fullAdder fa3_33 (.a(c2_18[12]) , .b(c2_18[11]) , .cin(c2_18[10]) , .s(c3_18[13]) , .c(c3_19[17]) ) ;

//idx19
fullAdder fa3_34 (.a(c2_19[19]) , .b(c2_19[18]) , .cin(c2_19[17]) , .s(c3_19[16]) , .c(c3_20[20]) ) ;
fullAdder fa3_35 (.a(c2_19[16]) , .b(c2_19[15]) , .cin(c2_19[14]) , .s(c3_19[15]) , .c(c3_20[19]) ) ;
fullAdder fa3_36 (.a(c2_19[13]) , .b(c2_19[12]) , .cin(c2_19[11]) , .s(c3_19[14]) , .c(c3_20[18]) ) ;

//idx20
fullAdder fa3_37 (.a(c2_20[20]) , .b(c2_20[19]) , .cin(c2_20[18]) , .s(c3_20[17]) , .c(c3_21[21]) ) ;
fullAdder fa3_38 (.a(c2_20[17]) , .b(c2_20[16]) , .cin(c2_20[15]) , .s(c3_20[16]) , .c(c3_21[20]) ) ;
fullAdder fa3_39 (.a(c2_20[14]) , .b(c2_20[13]) , .cin(c2_20[12]) , .s(c3_20[15]) , .c(c3_21[19]) ) ;

//idx21
fullAdder fa3_40 (.a(c2_21[21]) , .b(c2_21[20]) , .cin(c2_21[19]) , .s(c3_21[18]) , .c(c3_22[22]) ) ;
fullAdder fa3_41 (.a(c2_21[18]) , .b(c2_21[17]) , .cin(c2_21[16]) , .s(c3_21[17]) , .c(c3_22[21]) ) ;
fullAdder fa3_42 (.a(c2_21[15]) , .b(c2_21[14]) , .cin(c2_21[13]) , .s(c3_21[16]) , .c(c3_22[20]) ) ;

//idx22
fullAdder fa3_43 (.a(c2_22[22]) , .b(c2_22[21]) , .cin(c2_22[20]) , .s(c3_22[19]) , .c(c3_23[23]) ) ;
fullAdder fa3_44 (.a(c2_22[19]) , .b(c2_22[18]) , .cin(c2_22[17]) , .s(c3_22[18]) , .c(c3_23[22]) ) ;
fullAdder fa3_45 (.a(c2_22[16]) , .b(c2_22[15]) , .cin(c2_22[14]) , .s(c3_22[17]) , .c(c3_23[21]) ) ;

//idx23
fullAdder fa3_46 (.a(c2_23[23]) , .b(c2_23[22]) , .cin(c2_23[21]) , .s(c3_23[20]) , .c(c3_24[24]) ) ;
fullAdder fa3_47 (.a(c2_23[20]) , .b(c2_23[19]) , .cin(c2_23[18]) , .s(c3_23[19]) , .c(c3_24[23]) ) ;
fullAdder fa3_48 (.a(c2_23[17]) , .b(c2_23[16]) , .cin(c2_23[15]) , .s(c3_23[18]) , .c(c3_24[22]) ) ;

//idx24
fullAdder fa3_49 (.a(c2_24[24]) , .b(c2_24[23]) , .cin(c2_24[22]) , .s(c3_24[21]) , .c(c3_25[25]) ) ;
fullAdder fa3_50 (.a(c2_24[21]) , .b(c2_24[20]) , .cin(c2_24[19]) , .s(c3_24[20]) , .c(c3_25[24]) ) ;
assign c3_24[19]=c2_24[18];

//idx25
fullAdder fa3_51 (.a(c2_25[25]) , .b(c2_25[24]) , .cin(c2_25[23]) , .s(c3_25[23]) , .c(c3_26[26]) ) ;
assign c3_25[22:20]=c2_25[22:20];
assign c3_26[25:21]=c2_26[26:22]; assign c3_27 = c2_27; assign c3_28 = c2_28; assign c3_29 = c2_29; assign c3_30 = c2_30;


//stage4

wire  c4_0 ; wire [1:0] c4_1 ; wire [2:0] c4_2 ; wire [3:0] c4_3 ; wire [4:1] c4_4 ; wire [5:2] c4_5 ; wire [6:3] c4_6 ; wire [7:4] c4_7 ;
wire [8:5] c4_8 ; wire [9:6] c4_9 ; wire [10:7] c4_10 ; wire [11:8] c4_11 ; wire [12:9] c4_12 ; wire [13:10] c4_13 ; wire [14:11] c4_14 ; wire [15:12] c4_15 ; 
wire [16:13] c4_16 ; wire [17:14] c4_17 ; wire [18:15] c4_18 ; wire [19:16] c4_19 ; wire [20:17] c4_20 ; wire [21:18] c4_21 ; wire [22:19] c4_22 ;
wire [23:20] c4_23 ; wire [24:21] c4_24 ; wire [25:22] c4_25 ; wire [26:23] c4_26 ; wire [27:24] c4_27 ; wire [28:25] c4_28 ; wire [29:28] c4_29 ; wire c4_30;

assign c4_0 = c3_0 ; assign c4_1 = c3_1; assign c4_2 = c3_2 ; assign c4_3 = c3_3; 
//idx4
halfAdder ha4_1 (.a(c3_4[4]) , .b(c3_4[3]) , .s(c4_4[4]) , .c(c4_5[5]) ) ;
assign c4_4[3:1] = c3_4[2:0];

//idx5
fullAdder fa4_1 (.a(c3_5[5]) , .b(c3_5[4]) , .cin(c3_5[3]) , .s(c4_5[4]) , .c(c4_6[6]) ) ;
halfAdder ha4_2 (.a(c3_5[2]) , .b(c3_5[1]) , .s(c4_5[3]) , .c(c4_6[5]) ) ;
assign c4_5[2] = c3_5[0];

//idx6
fullAdder fa4_2 (.a(c3_6[6]) , .b(c3_6[5]) , .cin(c3_6[4]) , .s(c4_6[4]) , .c(c4_7[7]) ) ;
fullAdder fa4_3 (.a(c3_6[3]) , .b(c3_6[2]) , .cin(c3_6[1]) , .s(c4_6[3]) , .c(c4_7[6]) ) ;

//idx7
fullAdder fa4_4 (.a(c3_7[7]) , .b(c3_7[6]) , .cin(c3_7[5]) , .s(c4_7[5]) , .c(c4_8[8]) ) ;
fullAdder fa4_5 (.a(c3_7[4]) , .b(c3_7[3]) , .cin(c3_7[2]) , .s(c4_7[4]) , .c(c4_8[7]) ) ;
//idx8
fullAdder fa4_6 (.a(c3_8[8]) , .b(c3_8[7]) , .cin(c3_8[6]) , .s(c4_8[6]) , .c(c4_9[9]) ) ;
fullAdder fa4_7 (.a(c3_8[5]) , .b(c3_8[4]) , .cin(c3_8[3]) , .s(c4_8[5]) , .c(c4_9[8]) ) ;
//idx9
fullAdder fa4_8 (.a(c3_9[9]) , .b(c3_9[8]) , .cin(c3_9[7]) , .s(c4_9[7]) , .c(c4_10[10]) ) ;
fullAdder fa4_9 (.a(c3_9[6]) , .b(c3_9[5]) , .cin(c3_9[4]) , .s(c4_9[6]) , .c(c4_10[9]) ) ;

//idx10
fullAdder fa4_10 (.a(c3_10[10]) , .b(c3_10[9]) , .cin(c3_10[8]) , .s(c4_10[8]) , .c(c4_11[11]) ) ;
fullAdder fa4_11 (.a(c3_10[7]) , .b(c3_10[6]) , .cin(c3_10[5]) , .s(c4_10[7]) , .c(c4_11[10]) ) ;

//idx11
fullAdder fa4_12 (.a(c3_11[11]) , .b(c3_11[10]) , .cin(c3_11[9]) , .s(c4_11[9]) , .c(c4_12[12]) ) ;
fullAdder fa4_13 (.a(c3_11[8]) , .b(c3_11[7]) , .cin(c3_11[6]) , .s(c4_11[8]) , .c(c4_12[11]) ) ;

//idx12
fullAdder fa4_14 (.a(c3_12[12]) , .b(c3_12[11]) , .cin(c3_12[10]) , .s(c4_12[10]) , .c(c4_13[13]) ) ;
fullAdder fa4_15 (.a(c3_12[9]) , .b(c3_12[8]) , .cin(c3_12[7]) , .s(c4_12[9]) , .c(c4_13[12]) ) ;

//idx13
fullAdder fa4_16 (.a(c3_13[13]) , .b(c3_13[12]) , .cin(c3_13[11]) , .s(c4_13[11]) , .c(c4_14[14]) ) ;
fullAdder fa4_17 (.a(c3_13[10]) , .b(c3_13[9]) , .cin(c3_13[8]) , .s(c4_13[10]) , .c(c4_14[13]) ) ;

//idx14
fullAdder fa4_18 (.a(c3_14[14]) , .b(c3_14[13]) , .cin(c3_14[12]) , .s(c4_14[12]) , .c(c4_15[15]) ) ;
fullAdder fa4_19 (.a(c3_14[11]) , .b(c3_14[10]) , .cin(c3_14[9]) , .s(c4_14[11]) , .c(c4_15[14]) ) ;

//idx15
fullAdder fa4_20 (.a(c3_15[15]) , .b(c3_15[14]) , .cin(c3_15[13]) , .s(c4_15[13]) , .c(c4_16[16]) ) ;
fullAdder fa4_21 (.a(c3_15[12]) , .b(c3_15[11]) , .cin(c3_15[10]) , .s(c4_15[12]) , .c(c4_16[15]) ) ;

//idx16
fullAdder fa4_22 (.a(c3_16[16]) , .b(c3_16[15]) , .cin(c3_16[14]) , .s(c4_16[14]) , .c(c4_17[17]) ) ;
fullAdder fa4_23 (.a(c3_16[13]) , .b(c3_16[12]) , .cin(c3_16[11]) , .s(c4_16[13]) , .c(c4_17[16]) ) ;

//idx17
fullAdder fa4_24 (.a(c3_17[17]) , .b(c3_17[16]) , .cin(c3_17[15]) , .s(c4_17[15]) , .c(c4_18[18]) ) ;
fullAdder fa4_25 (.a(c3_17[14]) , .b(c3_17[13]) , .cin(c3_17[12]) , .s(c4_17[14]) , .c(c4_18[17]) ) ;

//idx18
fullAdder fa4_26 (.a(c3_18[18]) , .b(c3_18[17]) , .cin(c3_18[16]) , .s(c4_18[16]) , .c(c4_19[19]) ) ;
fullAdder fa4_27 (.a(c3_18[15]) , .b(c3_18[14]) , .cin(c3_18[13]) , .s(c4_18[15]) , .c(c4_19[18]) ) ;

//idx19
fullAdder fa4_28 (.a(c3_19[19]) , .b(c3_19[18]) , .cin(c3_19[17]) , .s(c4_19[17]) , .c(c4_20[20]) ) ;
fullAdder fa4_29 (.a(c3_19[16]) , .b(c3_19[15]) , .cin(c3_19[14]) , .s(c4_19[16]) , .c(c4_20[19]) ) ;

//idx20
fullAdder fa4_30 (.a(c3_20[20]) , .b(c3_20[19]) , .cin(c3_20[18]) , .s(c4_20[18]) , .c(c4_21[21]) ) ;
fullAdder fa4_31 (.a(c3_20[17]) , .b(c3_20[16]) , .cin(c3_20[15]) , .s(c4_20[17]) , .c(c4_21[20]) ) ;

//idx21
fullAdder fa4_32 (.a(c3_21[21]) , .b(c3_21[20]) , .cin(c3_21[19]) , .s(c4_21[19]) , .c(c4_22[22]) ) ;
fullAdder fa4_33 (.a(c3_21[18]) , .b(c3_21[17]) , .cin(c3_21[16]) , .s(c4_21[18]) , .c(c4_22[21]) ) ;

//idx22
fullAdder fa4_34 (.a(c3_22[22]) , .b(c3_22[21]) , .cin(c3_22[20]) , .s(c4_22[20]) , .c(c4_23[23]) ) ;
fullAdder fa4_35 (.a(c3_22[19]) , .b(c3_22[18]) , .cin(c3_22[17]) , .s(c4_22[19]) , .c(c4_23[22]) ) ;

//idx23
fullAdder fa4_36 (.a(c3_23[23]) , .b(c3_23[22]) , .cin(c3_23[21]) , .s(c4_23[21]) , .c(c4_24[24]) ) ;
fullAdder fa4_37 (.a(c3_23[20]) , .b(c3_23[19]) , .cin(c3_23[18]) , .s(c4_23[20]) , .c(c4_24[23]) ) ;

//idx24
fullAdder fa4_38 (.a(c3_24[24]) , .b(c3_24[23]) , .cin(c3_24[22]) , .s(c4_24[22]) , .c(c4_25[25]) ) ;
fullAdder fa4_39 (.a(c3_24[21]) , .b(c3_24[20]) , .cin(c3_24[19]) , .s(c4_24[21]) , .c(c4_25[24]) ) ;

//idx25
fullAdder fa4_40 (.a(c3_25[25]) , .b(c3_25[24]) , .cin(c3_25[23]) , .s(c4_25[23]) , .c(c4_26[26]) ) ;
fullAdder fa4_41 (.a(c3_25[22]) , .b(c3_25[21]) , .cin(c3_25[20]) , .s(c4_25[22]) , .c(c4_26[25]) ) ;

//idx26
fullAdder fa4_42 (.a(c3_26[26]) , .b(c3_26[25]) , .cin(c3_26[24]) , .s(c4_26[24]) , .c(c4_27[27]) ) ;
fullAdder fa4_43 (.a(c3_26[23]) , .b(c3_26[22]) , .cin(c3_26[21]) , .s(c4_26[23]) , .c(c4_27[26]) ) ;

//idx27
fullAdder fa4_44 (.a(c3_27[27]) , .b(c3_27[26]) , .cin(c3_27[25]) , .s(c4_27[25]) , .c(c4_28[28]) ) ;
assign c4_27[24]=c3_27[24];
assign c4_28[27:25]=c3_28[28:26] ; assign c4_29=c3_29; assign c4_30=c3_30 ;

//stage 5

wire  c5_0 ; wire [1:0] c5_1 ; wire [2:0] c5_2 ; wire [3:1] c5_3 ; wire [4:2] c5_4 ; wire [5:3] c5_5 ; wire [6:4] c5_6 ;wire [7:5] c5_7 ;wire [8:6] c5_8 ;
wire [9:7] c5_9 ;wire [10:8] c5_10 ;wire [11:9] c5_11 ;wire [12:10] c5_12 ;wire [13:11] c5_13 ;wire [14:12] c5_14 ;wire [15:13] c5_15 ;wire [16:14] c5_16 ;
wire [17:15] c5_17 ;wire [18:16] c5_18 ;wire [19:17] c5_19 ;wire [20:18] c5_20 ;wire [21:19] c5_21 ;wire [22:20] c5_22 ;
wire [23:21] c5_23 ;wire [24:22] c5_24 ;wire [25:23] c5_25 ;wire [26:24] c5_26 ;wire [27:25] c5_27 ;wire [28:26] c5_28 ;wire [29:27] c5_29 ; wire c5_30 ;
assign c5_0 = c4_0 ; assign c5_1=c4_1; assign c5_2 = c4_2;

halfAdder ha5_1 (.a(c4_3[3]) , .b(c4_3[2])  , .s(c5_3[3]) , .c(c5_4[4]) ) ;
assign c5_3[2:1]=c4_3[1:0];

fullAdder fa5_1 (.a(c4_4[4]) , .b(c4_4[3]) , .cin(c4_4[2]) , .s(c5_4[3]) , .c(c5_5[5]) ) ;
assign c5_4[2]=c4_4[1];

fullAdder fa5_2 (.a(c4_5[5]) , .b(c4_5[4]) , .cin(c4_5[3]) , .s(c5_5[4]) , .c(c5_6[6]) ) ;
assign c5_5[3]=c4_5[2];

fullAdder fa5_3 (.a(c4_6[6]) , .b(c4_6[5]) , .cin(c4_6[4]) , .s(c5_6[5]) , .c(c5_7[7]) ) ;
assign c5_6[4]=c4_6[3];

fullAdder fa5_4 (.a(c4_7[7]) , .b(c4_7[6]) , .cin(c4_7[5]) , .s(c5_7[6]) , .c(c5_8[8]) ) ;
assign c5_7[5] = c4_7[4];

fullAdder fa5_5 (.a(c4_8[8]) , .b(c4_8[7]) , .cin(c4_8[6]) , .s(c5_8[7]) , .c(c5_9[9]) ) ;
assign c5_8[6] = c4_8[5];

fullAdder fa5_6 (.a(c4_9[9]) , .b(c4_9[8]) , .cin(c4_9[7]) , .s(c5_9[8]) , .c(c5_10[10]) ) ;
assign c5_9[7] = c4_9[6];

fullAdder fa5_7 (.a(c4_10[10]) , .b(c4_10[9]) , .cin(c4_10[8]) , .s(c5_10[9]) , .c(c5_11[11]) ) ;
assign c5_10[8] = c4_10[7];

fullAdder fa5_8 (.a(c4_11[11]) , .b(c4_11[10]) , .cin(c4_11[9]) , .s(c5_11[10]) , .c(c5_12[12]) ) ;
assign c5_11[9] = c4_11[8];

fullAdder fa5_9 (.a(c4_12[12]) , .b(c4_12[11]) , .cin(c4_12[10]) , .s(c5_12[11]) , .c(c5_13[13]) ) ;
assign c5_12[10] = c4_12[9];

fullAdder fa5_10 (.a(c4_13[13]) , .b(c4_13[12]) , .cin(c4_13[11]) , .s(c5_13[12]) , .c(c5_14[14]) ) ;
assign c5_13[11] = c4_13[10];

fullAdder fa5_11 (.a(c4_14[14]) , .b(c4_14[13]) , .cin(c4_14[12]) , .s(c5_14[13]) , .c(c5_15[15]) ) ;
assign c5_14[12] = c4_14[11];

fullAdder fa5_12 (.a(c4_15[15]) , .b(c4_15[14]) , .cin(c4_15[13]) , .s(c5_15[14]) , .c(c5_16[16]) ) ;
assign c5_15[13] = c4_15[12];

fullAdder fa5_13 (.a(c4_16[16]) , .b(c4_16[15]) , .cin(c4_16[14]) , .s(c5_16[15]) , .c(c5_17[17]) ) ;
assign c5_16[14] = c4_16[13];

fullAdder fa5_14 (.a(c4_17[17]) , .b(c4_17[16]) , .cin(c4_17[15]) , .s(c5_17[16]) , .c(c5_18[18]) ) ;
assign c5_17[15] = c4_17[14];

fullAdder fa5_15 (.a(c4_18[18]) , .b(c4_18[17]) , .cin(c4_18[16]) , .s(c5_18[17]) , .c(c5_19[19]) ) ;
assign c5_18[16] = c4_18[15];

fullAdder fa5_16 (.a(c4_19[19]) , .b(c4_19[18]) , .cin(c4_19[17]) , .s(c5_19[18]) , .c(c5_20[20]) ) ;
assign c5_19[17] = c4_19[16];

fullAdder fa5_17 (.a(c4_20[20]) , .b(c4_20[19]) , .cin(c4_20[18]) , .s(c5_20[19]) , .c(c5_21[21]) ) ;
assign c5_20[18] = c4_20[17];

fullAdder fa5_18 (.a(c4_21[21]) , .b(c4_21[20]) , .cin(c4_21[19]) , .s(c5_21[20]) , .c(c5_22[22]) ) ;
assign c5_21[19] = c4_21[18];

fullAdder fa5_19 (.a(c4_22[22]) , .b(c4_22[21]) , .cin(c4_22[20]) , .s(c5_22[21]) , .c(c5_23[23]) ) ;
assign c5_22[20] = c4_22[19];

fullAdder fa5_20 (.a(c4_23[23]) , .b(c4_23[22]) , .cin(c4_23[21]) , .s(c5_23[22]) , .c(c5_24[24]) ) ;
assign c5_23[21] = c4_23[20];

fullAdder fa5_21 (.a(c4_24[24]) , .b(c4_24[23]) , .cin(c4_24[22]) , .s(c5_24[23]) , .c(c5_25[25]) ) ;
assign c5_24[22] = c4_24[21];

fullAdder fa5_22 (.a(c4_25[25]) , .b(c4_25[24]) , .cin(c4_25[23]) , .s(c5_25[24]) , .c(c5_26[26]) ) ;
assign c5_25[23] = c4_25[22];

fullAdder fa5_23 (.a(c4_26[26]) , .b(c4_26[25]) , .cin(c4_26[24]) , .s(c5_26[25]) , .c(c5_27[27]) ) ;
assign c5_26[24] = c4_26[23];

fullAdder fa5_24 (.a(c4_27[27]) , .b(c4_27[26]) , .cin(c4_27[25]) , .s(c5_27[26]) , .c(c5_28[28]) ) ;
assign c5_27[25] = c4_27[24];

fullAdder fa5_25 (.a(c4_28[28]) , .b(c4_28[27]) , .cin(c4_28[26]) , .s(c5_28[27]) , .c(c5_29[29]) ) ;
assign c5_28[26] = c4_28[25]; assign c5_29[28:27]=c4_29[29:28] ; assign c5_30=c4_30  ;

//stage 6
wire  c6_0 ; wire [1:0] c6_1 ; wire [2:1] c6_2 ; wire [3:2] c6_3 ; wire [4:3] c6_4 ; wire [5:4] c6_5 ; wire [6:5] c6_6 ;
wire [7:6] c6_7 ;wire [8:7] c6_8 ;wire [9:8] c6_9 ; wire [10:9] c6_10 ; wire [11:10] c6_11 ; wire [12:11] c6_12 ;
wire [13:12] c6_13 ; wire [14:13] c6_14 ; wire [15:14] c6_15 ; wire [16:15] c6_16 ; wire [17:16] c6_17 ; wire [18:17] c6_18 ; wire [19:18] c6_19 ;
wire [20:19] c6_20 ; wire [21:20] c6_21 ; wire [22:21] c6_22 ; wire [23:22] c6_23 ; wire [24:23] c6_24 ; wire [25:24] c6_25 ; wire [26:25] c6_26 ;
wire [27:26] c6_27 ; wire [28:27] c6_28 ; wire [29:28] c6_29 ; wire [30:29] c6_30 ;

assign c6_0 = c5_0; assign c6_1 = c5_1 ;
halfAdder ha6_1 (.a(c5_2[2]) , .b(c5_2[1])  , .s(c6_2[2]) , .c(c6_3[3]) ) ;
assign c6_2[1]=c5_2[0];

fullAdder fa6_1 (.a(c5_3[3]) , .b(c5_3[2]) , .cin(c5_3[1]) , .s(c6_3[2]) , .c(c6_4[4]) ) ;
fullAdder fa6_2 (.a(c5_4[4]) , .b(c5_4[3]) , .cin(c5_4[2]) , .s(c6_4[3]) , .c(c6_5[5]) ) ;
fullAdder fa6_3 (.a(c5_5[5]) , .b(c5_5[4]) , .cin(c5_5[3]) , .s(c6_5[4]) , .c(c6_6[6]) ) ;
fullAdder fa6_4 (.a(c5_6[6]) , .b(c5_6[5]) , .cin(c5_6[4]) , .s(c6_6[5]) , .c(c6_7[7]) ) ;
fullAdder fa6_5 (.a(c5_7[7]) , .b(c5_7[6]) , .cin(c5_7[5]) , .s(c6_7[6]) , .c(c6_8[8]) ) ;
fullAdder fa6_6 (.a(c5_8[8]) , .b(c5_8[7]) , .cin(c5_8[6]) , .s(c6_8[7]) , .c(c6_9[9]) ) ;
fullAdder fa6_7 (.a(c5_9[9]) , .b(c5_9[8]) , .cin(c5_9[7]) , .s(c6_9[8]) , .c(c6_10[10]) ) ;
fullAdder fa6_8 (.a(c5_10[10]) , .b(c5_10[9]) , .cin(c5_10[8]) , .s(c6_10[9]) , .c(c6_11[11]) ) ;
fullAdder fa6_9 (.a(c5_11[11]) , .b(c5_11[10]) , .cin(c5_11[9]) , .s(c6_11[10]) , .c(c6_12[12]) ) ;
fullAdder fa6_10 (.a(c5_12[12]) , .b(c5_12[11]) , .cin(c5_12[10]) , .s(c6_12[11]) , .c(c6_13[13]) ) ;
fullAdder fa6_11 (.a(c5_13[13]) , .b(c5_13[12]) , .cin(c5_13[11]) , .s(c6_13[12]) , .c(c6_14[14]) ) ;
fullAdder fa6_12 (.a(c5_14[14]) , .b(c5_14[13]) , .cin(c5_14[12]) , .s(c6_14[13]) , .c(c6_15[15]) ) ;
fullAdder fa6_13 (.a(c5_15[15]) , .b(c5_15[14]) , .cin(c5_15[13]) , .s(c6_15[14]) , .c(c6_16[16]) ) ;
fullAdder fa6_14 (.a(c5_16[16]) , .b(c5_16[15]) , .cin(c5_16[14]) , .s(c6_16[15]) , .c(c6_17[17]) ) ;
fullAdder fa6_15 (.a(c5_17[17]) , .b(c5_17[16]) , .cin(c5_17[15]) , .s(c6_17[16]) , .c(c6_18[18]) ) ;
fullAdder fa6_16 (.a(c5_18[18]) , .b(c5_18[17]) , .cin(c5_18[16]) , .s(c6_18[17]) , .c(c6_19[19]) ) ;
fullAdder fa6_17 (.a(c5_19[19]) , .b(c5_19[18]) , .cin(c5_19[17]) , .s(c6_19[18]) , .c(c6_20[20]) ) ;
fullAdder fa6_18 (.a(c5_20[20]) , .b(c5_20[19]) , .cin(c5_20[18]) , .s(c6_20[19]) , .c(c6_21[21]) ) ;
fullAdder fa6_19 (.a(c5_21[21]) , .b(c5_21[20]) , .cin(c5_21[19]) , .s(c6_21[20]) , .c(c6_22[22]) ) ;
fullAdder fa6_20 (.a(c5_22[22]) , .b(c5_22[21]) , .cin(c5_22[20]) , .s(c6_22[21]) , .c(c6_23[23]) ) ;
fullAdder fa6_21 (.a(c5_23[23]) , .b(c5_23[22]) , .cin(c5_23[21]) , .s(c6_23[22]) , .c(c6_24[24]) ) ;
fullAdder fa6_22 (.a(c5_24[24]) , .b(c5_24[23]) , .cin(c5_24[22]) , .s(c6_24[23]) , .c(c6_25[25]) ) ;
fullAdder fa6_23 (.a(c5_25[25]) , .b(c5_25[24]) , .cin(c5_25[23]) , .s(c6_25[24]) , .c(c6_26[26]) ) ;
fullAdder fa6_24 (.a(c5_26[26]) , .b(c5_26[25]) , .cin(c5_26[24]) , .s(c6_26[25]) , .c(c6_27[27]) ) ;
fullAdder fa6_25 (.a(c5_27[27]) , .b(c5_27[26]) , .cin(c5_27[25]) , .s(c6_27[26]) , .c(c6_28[28]) ) ;
fullAdder fa6_26 (.a(c5_28[28]) , .b(c5_28[27]) , .cin(c5_28[26]) , .s(c6_28[27]) , .c(c6_29[29]) ) ;
fullAdder fa6_27 (.a(c5_29[29]) , .b(c5_29[28]) , .cin(c5_29[27]) , .s(c6_29[28]) , .c(c6_30[30]) ) ;
assign c6_30[29]=c5_30 ;

wire [31:0] r1 ;
wire [31:0] r2 ;
assign r1[0]=c6_0; assign r2[0]= 0 ;
assign r1[31]=0; assign r2[31]= 0 ;
assign r1[30:1] = {c6_30[30], c6_29[29], c6_28[28], c6_27[27], c6_26[26], c6_25[25], c6_24[24], c6_23[23], c6_22[22], c6_21[21], c6_20[20], c6_19[19], c6_18[18], c6_17[17], c6_16[16], c6_15[15], c6_14[14], c6_13[13], c6_12[12], c6_11[11], c6_10[10], c6_9[9], c6_8[8], c6_7[7], c6_6[6], c6_5[5], c6_4[4], c6_3[3], c6_2[2], c6_1[1]};
assign r2[30:1] = {c6_30[29], c6_29[28], c6_28[27], c6_27[26], c6_26[25], c6_25[24], c6_24[23], c6_23[22], c6_22[21], c6_21[20], c6_20[19], c6_19[18], c6_18[17], c6_17[16], c6_16[15], c6_15[14], c6_14[13], c6_13[12], c6_12[11], c6_11[10], c6_10[9], c6_9[8], c6_8[7], c6_7[6], c6_6[5], c6_5[4], c6_4[3], c6_3[2], c6_2[1], c6_1[0]};

//assign y = r1+r2 ;

brentkung bk(.a(r1),.b(r2),.cin(0),.sum(y[30:0]),.cout(y[31]));

//always @(*) begin
//  $display("Stage0:\n c0_0= %b | c0_1= %b | c0_2= %b | c0_3= %b | c0_4= %b | c0_5= %b | c0_6= %b | c0_7= %b\n \
//            c0_8= %b | c0_9= %b | c0_10= %b | c0_11= %b | c0_12= %b | c0_13= %b | c0_14= %b | c0_15= %b\n \
//            c0_16= %b | c0_17= %b | c0_18= %b | c0_19= %b | c0_20= %b | c0_21= %b | c0_22= %b | c0_23= %b\n \
//            c0_24= %b | c0_25= %b | c0_26= %b | c0_27= %b | c0_28= %b | c0_29= %b | c0_30= %b\n\n \
//Stage1:\n c1_0= %b | c1_1= %b | c1_2= %b | c1_3= %b | c1_4= %b | c1_5= %b | c1_6= %b | c1_7= %b\n \
//            c1_8= %b | c1_9= %b | c1_10= %b | c1_11= %b | c1_12= %b | c1_13= %b | c1_14= %b | c1_15= %b\n \
//            c1_16= %b | c1_17= %b | c1_18= %b | c1_19= %b | c1_20= %b | c1_21= %b | c1_22= %b | c1_23= %b\n \
//            c1_24= %b | c1_25= %b | c1_26= %b | c1_27= %b | c1_28= %b | c1_29= %b | c1_30= %b\n\n \
//Stage2:\n c2_0= %b | c2_1= %b | c2_2= %b | c2_3= %b | c2_4= %b | c2_5= %b | c2_6= %b | c2_7= %b\n \
//            c2_8= %b | c2_9= %b | c2_10= %b | c2_11= %b | c2_12= %b | c2_13= %b | c2_14= %b | c2_15= %b\n \
//            c2_16= %b | c2_17= %b | c2_18= %b | c2_19= %b | c2_20= %b | c2_21= %b | c2_22= %b | c2_23= %b\n \
//            c2_24= %b | c2_25= %b | c2_26= %b | c2_27= %b | c2_28= %b | c2_29= %b | c2_30= %b\n\n \
//Stage3:\n c3_0= %b | c3_1= %b | c3_2= %b | c3_3= %b | c3_4= %b | c3_5= %b | c3_6= %b | c3_7= %b\n \
//            c3_8= %b | c3_9= %b | c3_10= %b | c3_11= %b | c3_12= %b | c3_13= %b | c3_14= %b | c3_15= %b\n \
//            c3_16= %b | c3_17= %b | c3_18= %b | c3_19= %b | c3_20= %b | c3_21= %b | c3_22= %b | c3_23= %b\n \
//            c3_24= %b | c3_25= %b | c3_26= %b | c3_27= %b | c3_28= %b | c3_29= %b | c3_30= %b\n\n \
//Stage4:\n c4_0= %b | c4_1= %b | c4_2= %b | c4_3= %b | c4_4= %b | c4_5= %b | c4_6= %b | c4_7= %b\n \
//            c4_8= %b | c4_9= %b | c4_10= %b | c4_11= %b | c4_12= %b | c4_13= %b | c4_14= %b | c4_15= %b\n \
//            c4_16= %b | c4_17= %b | c4_18= %b | c4_19= %b | c4_20= %b | c4_21= %b | c4_22= %b | c4_23= %b\n \
//            c4_24= %b | c4_25= %b | c4_26= %b | c4_27= %b | c4_28= %b | c4_29= %b | c4_30= %b\n\n \
//Stage5:\n c5_0= %b | c5_1= %b | c5_2= %b | c5_3= %b | c5_4= %b | c5_5= %b | c5_6= %b | c5_7= %b\n \
//            c5_8= %b | c5_9= %b | c5_10= %b | c5_11= %b | c5_12= %b | c5_13= %b | c5_14= %b | c5_15= %b\n \
//            c5_16= %b | c5_17= %b | c5_18= %b | c5_19= %b | c5_20= %b | c5_21= %b | c5_22= %b | c5_23= %b\n \
//            c5_24= %b | c5_25= %b | c5_26= %b | c5_27= %b | c5_28= %b | c5_29= %b | c5_30= %b\n\n \
//Stage6:\n c6_0= %b | c6_1= %b | c6_2= %b | c6_3= %b | c6_4= %b | c6_5= %b | c6_6= %b | c6_7= %b\n \
//            c6_8= %b | c6_9= %b | c6_10= %b | c6_11= %b | c6_12= %b | c6_13= %b | c6_14= %b | c6_15= %b\n \
//            c6_16= %b | c6_17= %b | c6_18= %b | c6_19= %b | c6_20= %b | c6_21= %b | c6_22= %b | c6_23= %b\n \
//            c6_24= %b | c6_25= %b | c6_26= %b | c6_27= %b | c6_28= %b | c6_29= %b | c6_30= %b", 
//            c0_0, c0_1, c0_2, c0_3, c0_4, c0_5, c0_6, c0_7, 
//            c0_8, c0_9, c0_10, c0_11, c0_12, c0_13, c0_14, c0_15, 
//            c0_16, c0_17, c0_18, c0_19, c0_20, c0_21, c0_22, c0_23, 
//            c0_24, c0_25, c0_26, c0_27, c0_28, c0_29, c0_30, 
//            c1_0, c1_1, c1_2, c1_3, c1_4, c1_5, c1_6, c1_7, 
//            c1_8, c1_9, c1_10, c1_11, c1_12, c1_13, c1_14, c1_15, 
//            c1_16, c1_17, c1_18, c1_19, c1_20, c1_21, c1_22, c1_23, 
//            c1_24, c1_25, c1_26, c1_27, c1_28, c1_29, c1_30, 
//            c2_0, c2_1, c2_2, c2_3, c2_4, c2_5, c2_6, c2_7, 
//            c2_8, c2_9, c2_10, c2_11, c2_12, c2_13, c2_14, c2_15, 
//            c2_16, c2_17, c2_18, c2_19, c2_20, c2_21, c2_22, c2_23, 
//            c2_24, c2_25, c2_26, c2_27, c2_28, c2_29, c2_30, 
//            c3_0, c3_1, c3_2, c3_3, c3_4, c3_5, c3_6, c3_7, 
//            c3_8, c3_9, c3_10, c3_11, c3_12, c3_13, c3_14, c3_15, 
//            c3_16, c3_17, c3_18, c3_19, c3_20, c3_21, c3_22, c3_23, 
//            c3_24, c3_25, c3_26, c3_27, c3_28, c3_29, c3_30, 
//            c4_0, c4_1, c4_2, c4_3, c4_4, c4_5, c4_6, c4_7, 
//            c4_8, c4_9, c4_10, c4_11, c4_12, c4_13, c4_14, c4_15, 
//            c4_16, c4_17, c4_18, c4_19, c4_20, c4_21, c4_22, c4_23, 
//            c4_24, c4_25, c4_26, c4_27, c4_28, c4_29, c4_30, 
//            c5_0, c5_1, c5_2, c5_3, c5_4, c5_5, c5_6, c5_7, 
//            c5_8, c5_9, c5_10, c5_11, c5_12, c5_13, c5_14, c5_15, 
//            c5_16, c5_17, c5_18, c5_19, c5_20, c5_21, c5_22, c5_23, 
//            c5_24, c5_25, c5_26, c5_27, c5_28, c5_29, c5_30, 
//            c6_0, c6_1, c6_2, c6_3, c6_4, c6_5, c6_6, c6_7, 
//            c6_8, c6_9, c6_10, c6_11, c6_12, c6_13, c6_14, c6_15, 
//            c6_16, c6_17, c6_18, c6_19, c6_20, c6_21, c6_22, c6_23, 
//            c6_24, c6_25, c6_26, c6_27, c6_28, c6_29, c6_30);
            
                                                   
//$display("Stage7:\n r1= %b | r2= %b", r1, r2);       
//end




endmodule

